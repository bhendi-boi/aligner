`include "./rtl/cfs_synch.sv"
`include "./rtl/cfs_synch_fifo.sv"
`include "./rtl/cfs_rx_ctrl.sv"
`include "./rtl/cfs_ctrl.sv"
`include "./rtl/cfs_tx_ctrl.sv"
`include "./rtl/cfs_edge_detect.sv"
`include "./rtl/cfs_regs.sv"
`include "./rtl/cfs_aligner_core.sv"
`include "./rtl/cfs_aligner.sv"
